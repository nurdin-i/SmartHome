module SmartHome
(
	input clk,
	output led1
);


main MAIN(
	.clk(clk),
	.led1(led1)
);

endmodule